module encoder(
    input wire [9:0]Keypad,
    input wire Clk,
    input wire Enablen,
    output wire [3:0]D,
    output wire loadn,
    output wire pgt_1Hz
);
    //TODO encoder
endmodule