module timer(

);

endmodule;