module microwave(
    input wire keypad[9:0],
    input wire clk,
    input wire startn,
    input wire stopn,
    input wire clearn,
    input wire door_closed,
    input wire timer_done
);


endmodule